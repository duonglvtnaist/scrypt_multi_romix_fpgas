module salsa_20_8(
		input	wire 			clk,
		input	wire			init,
		input	wire			reset_n,
		input	wire 	[31:0]	x0,
		input	wire 	[31:0]	x1,
		input	wire 	[31:0]	x2,
		input	wire 	[31:0]	x3,
		input	wire 	[31:0]	x4,
		input	wire 	[31:0]	x5,
		input	wire 	[31:0]	x6,
		input	wire 	[31:0]	x7,
		input	wire 	[31:0]	x8,
		input	wire 	[31:0]	x9,
		input	wire 	[31:0]	x10,
		input	wire 	[31:0]	x11,
		input	wire 	[31:0]	x12,
		input	wire 	[31:0]	x13,
		input	wire 	[31:0]	x14,
		input	wire 	[31:0]	x15,		
		output	wire 	[31:0]	out0,
		output	wire 	[31:0]	out1,
		output	wire 	[31:0]	out2,
		output	wire 	[31:0]	out3,
		output	wire 	[31:0]	out4,
		output	wire 	[31:0]	out5,
		output	wire 	[31:0]	out6,
		output	wire 	[31:0]	out7,
		output	wire 	[31:0]	out8,
		output	wire 	[31:0]	out9,
		output	wire 	[31:0]	out10,
		output	wire 	[31:0]	out11,
		output	wire 	[31:0]	out12,
		output	wire 	[31:0]	out13,
		output	wire 	[31:0]	out14,
		output	wire 	[31:0]	out15,
		output 	wire			valid
);

		wire sel_in;
		// wire sel_order;
		wire write_temp;
	salsa_20_8_ct controller (
		.clk(clk),
		.init(init),
		.reset_n(reset_n),
		.write_temp(write_temp),
		.sel_in(sel_in),
		// .sel_order(sel_order),
		.valid(valid)
	);

	salsa_20_8_dp datapath (
		.clk(clk),
		.reset_n(reset_n),
		.write_temp(write_temp),
		.sel_in(sel_in),
		// .sel_order(sel_order),
		.x0		(x0	)		,
		.x1		(x1	)		,
		.x2		(x2	)		,
		.x3		(x3	)		,
		.x4		(x4	)		,
		.x5		(x5	)		,
		.x6		(x6	)		,
		.x7		(x7	)		,
		.x8		(x8	)		,
		.x9		(x9	)		,
		.x10	(x10)		,
		.x11	(x11)		,
		.x12	(x12)		,
		.x13	(x13)		,
		.x14	(x14)		,
		.x15	(x15)		,
		.out0	(out0)		,
		.out1	(out1)		,
		.out2	(out2)		,
		.out3	(out3)		,
		.out4	(out4)		,
		.out5	(out5)		,
		.out6	(out6)		,
		.out7	(out7)		,
		.out8	(out8)		,
		.out9	(out9)		,
		.out10	(out10)		,
		.out11	(out11)		,
		.out12	(out12)		,
		.out13	(out13)		,
		.out14	(out14)		,
		.out15	(out15)		,
		.valid	(valid)
	);
endmodule 

